module digit_sum_ar(
input logic [3:0] s_1, s_2,
output logic [4:0] sum);

	assign sum = s_1 + s_2;
	
endmodule